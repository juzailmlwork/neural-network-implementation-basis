module tb_top_module;
    reg clk;
    reg reset;
    reg rx;
    reg read_request;
    wire [3:0] digit_out;
    wire image_written;
    wire read_enable;
    wire NN_done;

    logic signed [7:0] data_8 [0:783] = '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 69, 100, 126, 127, 116, 53, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 109, 126, 126, 105, 103, 107, 126, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 126, 116, 44, 3, 0, 6, 101, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 126, 126, 91, 0, 0, 0, 0, 79, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 126, 126, 39, 0, 0, 0, 0, 31, 21, 110, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 127, 116, 19, 0, 0, 0, 0, 3, 106, 126, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 126, 126, 77, 15, 0, 0, 4, 77, 126, 126, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 126, 126, 113, 92, 66, 98, 126, 126, 126, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 59, 80, 118, 126, 126, 126, 113, 80, 122, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 0, 0, 30, 42, 37, 11, 8, 0, 89, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 64, 5, 0, 0, 0, 0, 0, 0, 0, 0, 115, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 126, 58, 0, 0, 0, 0, 0, 0, 0, 0, 78, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 126, 58, 0, 0, 0, 0, 0, 0, 0, 0, 58, 118, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 126, 31, 0, 0, 0, 0, 0, 0, 0, 0, 58, 117, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 126, 58, 0, 0, 0, 0, 0, 0, 0, 0, 110, 120, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 126, 122, 30, 0, 0, 0, 0, 0, 19, 116, 126, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 108, 126, 118, 64, 4, 0, 0, 15, 77, 126, 115, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 126, 126, 126, 98, 40, 92, 114, 126, 113, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 109, 126, 126, 126, 126, 126, 126, 59, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 27, 89, 73, 95, 58, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 };
    logic signed [7:0] data_4 [0:783] = '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 97, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 93, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98, 127, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 113, 120, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 126, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 127, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 127, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 127, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 127, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 126, 90, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 124, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 101, 127, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 115, 124, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 127, 127, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 115, 124, 0, 36, 76, 0, 0, 0, 0, 0, 0, 0, 0, 127, 116, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 115, 126, 120, 123, 28, 0, 0, 0, 0, 0, 0, 0, 0, 124, 127, 57, 3, 0, 5, 7, 7, 7, 7, 10, 55, 55, 37, 87, 124, 126, 88, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 122, 127, 102, 86, 115, 127, 127, 127, 127, 127, 127, 105, 88, 57, 86, 126, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 92, 105, 105, 88, 85, 105, 71, 57, 55, 9, 4, 0, 0, 67, 127, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 127, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 127, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 127, 98, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 105, 127, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 127, 105, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 110, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 };
    integer rx_index = 0;
    reg signed [7:0] data [0:783];

    top_module uut (
        .clk(clk),
        .reset(reset),
        .rx(rx),
        .read_request(read_request),
        .image_written(image_written),
        .read_enable(read_enable),
        .NN_done(NN_done),
        .digit_out(digit_out)
    );

    initial begin
        clk = 0;
        reset = 1;
        rx = 1; // Idle state
        read_request = 1;
        data = data_4;
        #20 reset = 0;

        // Transmit 784 bytes
        repeat (784) begin
                  rx = 0; // Start bit
                  #40 rx = data[rx_index][0]; 
                  #40 rx = data[rx_index][1]; 
                  #40 rx = data[rx_index][2];
                  #40 rx = data[rx_index][3];
                  #40 rx = data[rx_index][4];
                  #40 rx = data[rx_index][5];
                  #40 rx = data[rx_index][6];
                  #40 rx = data[rx_index][7];
                  #40 rx = 1; // Stop bit
                     $display("Index: %d, Data: %d", rx_index, data[rx_index]);
                    rx_index = rx_index + 1;
        end

        wait(NN_done);
//        #50reset=1;
//        #10 $finish;
//        data = data_8;
//        rx_index = 0;
//        #20 reset = 0;
        
//                // Transmit 784 bytes
//                repeat (784) begin
//                          rx = 0; // Start bit
//                          #40 rx = data[rx_index][0]; 
//                          #40 rx = data[rx_index][1]; 
//                          #40 rx = data[rx_index][2];
//                          #40 rx = data[rx_index][3];
//                          #40 rx = data[rx_index][4];
//                          #40 rx = data[rx_index][5];
//                          #40 rx = data[rx_index][6];
//                          #40 rx = data[rx_index][7];
//                          #40 rx = 1; // Stop bit
//                             $display("Index: %d, Data: %d", rx_index, data[rx_index]);
//                            rx_index = rx_index + 1;
//                end
//        wait(NN_done);
        #10 $finish;
    end

    always #5 clk = ~clk; 
endmodule
